module shiftreg
#(
    // * --------------------------------------------------------------------
    // * Parameters
    // * --------------------------------------------------------------------
    parameter                        NB_DATA   = 3
)
(
    // * --------------------------------------------------------------------
    // * Outputs
    // * --------------------------------------------------------------------
    output logic [ NB_DATA - 1 : 0 ] o_led          ,

    // * --------------------------------------------------------------------
    // * Inputs
    // * --------------------------------------------------------------------
    input  logic                     i_valid        ,

    // * --------------------------------------------------------------------
    // * Clock and reset
    // * --------------------------------------------------------------------
    input  logic                     i_reset        ,
    input  logic                     i_clock
) ;
    // * --------------------------------------------------------------------
    // * Internal logics
    // * --------------------------------------------------------------------
    logic        [ NB_DATA - 1 : 0 ] shift_register ;

    // * --------------------------------------------------------------------
    // * Shift register
    // * --------------------------------------------------------------------
    always_ff @(posedge i_clock)
    begin : proc_data_move
        if (i_reset)
            shift_register <= {{NB_DATA-1{1'b0}}, 1'b1};
        else if (i_valid)
            shift_register <= {shift_register[NB_DATA-2:0], shift_register[NB_DATA-1]};
    end

    // * --------------------------------------------------------------------
    // * Output assignment
    // * --------------------------------------------------------------------
    assign o_led = shift_register;
endmodule
